module lab3_top_tb();

reg [9:0] SW;
reg [3:0] KEY;
reg [3:0] states;

wire [6:0] HEX0, HEX1, HEX2, HEX3, HEX4, HEX5;
wire [9:0] LEDR;

lab3_top DUT(SW,KEY,HEX0,HEX1,HEX2,HEX3,HEX4,HEX5,LEDR);

initial begin
SW = 10'b0;
KEY = 4'b0;

#5;

SW = {6'b000000,4'b0001};
KEY[3] = 1'b1;

$display ("Output is %b and in state %b, expected %b and %b",HEX0,states,7'b0110000,4'b1000);

#5;

SW = {6'b000000,4'b0001};
KEY[3] = 1'b1;

$display ("Output is %b and in state %b, expected %b and %b",HEX0,states,7'b0110000,4'b1000);

#5;

SW = {6'b000000,4'b1111};
KEY[0] = 1'b1;


$display ("Output is %b and in state %b, expected %b and %b",HEX0,states,7'b1111111,4'b0000);

#5;
SW = {6'b000000,4'b1111};
KEY[3] = 1'b1;

$display ("Output is %b and in state %b, expected %b and %b",HEX0,states,7'b1111111,4'b0001);
$stop;
end
endmodule
