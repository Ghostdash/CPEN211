module lab5_top_tb;
  reg [3:0] KEY;
  reg [9:0] SW;
  wire [9:0] LEDR; 
  wire [6:0] HEX0, HEX1, HEX2, HEX3, HEX4, HEX5;
  reg CLOCK_50;
  reg [2:0] debug;

  lab5_top DUT(KEY,SW,LEDR,HEX0,HEX1,HEX2,HEX3,HEX4,HEX5,CLOCK_50);

//  initial forever begin
//    CLOCK_50 = 0; #5;
//    CLOCK_50 = 1; #5;
//  end

  initial begin
	SW = 10'b1001000010;     //42 hex
	CLOCK_50 = 0;
#1;
	SW[9] = 1'b0;
#1;
	SW = 10'b0000010001;     //write to r2
#3;
	CLOCK_50 = 1;
#5;
	CLOCK_50 = 0;
#5;
 	SW = 10'b0000100000;      //load in A
#5;
	CLOCK_50 = 1;
#5;
	CLOCK_50 = 0;
	SW = 10'b1000010011;     //13
#1;
	SW[9] = 1'b0;
#1;
	SW = 10'b0000010011;     //write to r1
#3;
	CLOCK_50 = 1;
#5;
	CLOCK_50 = 0;
	SW = 10'b0001000010;     //load in B
#5;
	CLOCK_50 = 1;
#5;
	CLOCK_50 =0 ;
	SW = 10'b0010000000;      //load C
#5;
	CLOCK_50 =1;
#5;
	CLOCK_50 = 0;
$display("Output is %b, expecting %b",HEX0,7'b0010010);   //5
$display("Output is %b, expecting %b",HEX1,7'b0010010);   //5
    $stop;
  end
endmodule
