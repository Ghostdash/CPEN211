module lab7_top(KEY,SW,LEDR,HEX0,HEX1,HEX2,HEX3,HEX4,HEX5);
input [3:0] KEY;
input [9:0] SW;
output [9:0] LEDR;
output [6:0] HEX0, HEX1, HEX2, HEX3, HEX4, HEX5;

wire Z, N, V;
wire [8:0] mem_addr;
wire [1:0] mem_cmd;
wire [7:0] write_address;
wire [15:0] dout,din;

wire [15:0] out_mem,out_hex;

wire write,enable,msel,mread,mwrite;
wire zero;

assign zero = 1'b0;                               //a 1 bit wire set to zero for msel equal comparator
assign write_address = mem_addr[7:0];

EqComp #1 MSEL (mem_addr[8],zero,msel);         //equal comparators
EqComp #2 MREAD (mem_cmd,2'b10,mread);
EqComp #2 MWRITE (mem_cmd,2'b11,mwrite);

assign write = mwrite & msel;

assign enable = mread & msel;
assign out_mem = enable ? dout:{16{1'bz}}; //tri state enabler


  cpu CPU( .clk   (~KEY[0]), // recall from Lab 4 that KEY0 is 1 when NOT pushed
         .reset (~KEY[1]), 
         .load  (~KEY[3]),
         .in (out_mem),
	 .mdata (out_mem),
         .out   (out_hex),
         .Z     (Z),
         .N     (N),
         .V     (V),
         .w     (LEDR[9]), 
	 .mem_addr (mem_addr), 
	 .mem_cmd(mem_cmd)
	 );

RAM MEM(~KEY[0],mem_addr[7:0],write_address,write,out_hex,dout);

assign HEX5[0] = ~Z;
assign HEX5[6] = ~N;
assign HEX5[3] = ~V;

sseg H0(out_hex[3:0],   HEX0);
sseg H1(out_hex[7:4],   HEX1);
sseg H2(out_hex[11:8],  HEX2);
sseg H3(out_hex[15:12], HEX3);
  
assign HEX4 = 7'b1111111;
assign {HEX5[2:1],HEX5[5:4]} = 4'b1111; // disabled
assign LEDR[8] = 1'b0;

endmodule


// To ensure Quartus uses the embedded MLAB memory blocks inside the Cyclone
// V on your DE1-SoC we follow the coding style from in Altera's Quartus II
// Handbook (QII5V1 2015.05.04) in Chapter 12, ?Recommended HDL Coding Style?
//
// 1. "Example 12-11: Verilog Single Clock Simple Dual-Port Synchronous RAM 
//     with Old Data Read-During-Write Behavior" 
// 2. "Example 12-29: Verilog HDL RAM Initialized with the readmemb Command"

module RAM(clk,read_address,write_address,write,din,dout);
  parameter data_width = 16; 
  parameter addr_width = 8;
  parameter filename = "data.txt";

  input clk;
  input [addr_width-1:0] read_address, write_address;
  input write;
  input [data_width-1:0] din;
  output [data_width-1:0] dout;
  reg [data_width-1:0] dout;

  reg [data_width-1:0] mem [2**addr_width-1:0];

  initial $readmemb(filename, mem);

  always @ (posedge clk) begin
    if (write)
      mem[write_address] <= din;
    dout <= mem[read_address]; // dout doesn't get din in this clock cycle 
                               // (this is due to Verilog non-blocking assignment "<=")
  end 
endmodule



module sseg(in,segs);
  input [3:0] in;
  output [6:0] segs;

  reg [6:0] segs;

  // NOTE: The code for sseg below is not complete: You can use your code from
  // Lab4 to fill this in or code from someone else's Lab4.  
  //
  // IMPORTANT:  If you *do* use someone else's Lab4 code for the seven
  // segment display you *need* to state the following three things in
  // a file README.txt that you submit with handin along with this code: 
  //
  //   1.  First and last name of student providing code
  //   2.  Student number of student providing code
  //   3.  Date and time that student provided you their code
  //
  // You must also (obviously!) have the other student's permission to use
  // their code.
  //
  // To do otherwise is considered plagiarism.
  //
  // One bit per segment. On the DE1-SoC a HEX segment is illuminated when
  // the input bit is 0. Bits 6543210 correspond to:
  //
  //    0000
  //   5    1
  //   5    1
  //    6666
  //   4    2
  //   4    2
  //    3333
  //
  // Decimal value | Hexadecimal symbol to render on (one) HEX display
  //             0 | 0
  //             1 | 1
  //             2 | 2
  //             3 | 3
  //             4 | 4
  //             5 | 5
  //             6 | 6
  //             7 | 7
  //             8 | 8
  //             9 | 9
  //            10 | A
  //            11 | b
  //            12 | C
  //            13 | d
  //            14 | E
  //            15 | F
always @(*)
  case(in)
	4'b0000: segs = 7'b1000000;  //0
	4'b0001: segs = 7'b1111001;  //1
	4'b0010: segs = 7'b0100100;  //2
	4'b0011: segs = 7'b0110000;  //3
	4'b0100: segs = 7'b0011001;  //4
	4'b0101: segs = 7'b0010010;  //5
	4'b0110: segs = 7'b0000010;
	4'b0111: segs = 7'b1111000;
	4'b1000: segs = 7'b0000000;
	4'b1001: segs = 7'b0010000;
	4'b1010: segs = 7'b0001000;
	4'b1011: segs = 7'b0000011;
	4'b1100: segs = 7'b1000110;
	4'b1101: segs = 7'b0100001;
	4'b1110: segs = 7'b0000110;
	4'b1111: segs = 7'b0001110;
  default: segs = 7'b1000000;   //output "0"
endcase
endmodule

module EqComp(a, b, eq) ;
  parameter k=8;
  input  [k-1:0] a,b;
  output eq;
  wire   eq;

  assign eq = (a==b) ;
endmodule

